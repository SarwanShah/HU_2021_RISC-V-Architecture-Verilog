module top
(
	

);


endmodule 